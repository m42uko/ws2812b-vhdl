-- ----------------------------------------------------------------------------
--                         WS2812B CONTROLLER FOR FPGAS                        
-- ----------------------------------------------------------------------------
-- ws2812b_gamma.vhd : Gamma correction RAM for the WS2812B LEDs.
--                   : Do note that this generates a (fairly large, async) LUT.
-- ----------------------------------------------------------------------------
-- Author          : Markus Koch <markus@notsyncing.net>
-- Contributors    : None 
-- Created on      : 2016/10/16
-- License         : Mozilla Public License (MPL) Version 2
-- ----------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity ws2812b_gamma is
	port(
		pixelData_in  : in  std_logic_vector(7 downto 0);
		pixelData_out : out std_logic_vector(7 downto 0)
	);
end entity ws2812b_gamma;

architecture RTL of ws2812b_gamma is
	type gamma_table_t is array (0 to 255) of std_logic_vector(7 downto 0);
	constant gamma_table : gamma_table_t := (
		0   => std_logic_vector(to_unsigned(0, 8)),
		1   => std_logic_vector(to_unsigned(0, 8)),
		2   => std_logic_vector(to_unsigned(0, 8)),
		3   => std_logic_vector(to_unsigned(0, 8)),
		4   => std_logic_vector(to_unsigned(0, 8)),
		5   => std_logic_vector(to_unsigned(0, 8)),
		6   => std_logic_vector(to_unsigned(0, 8)),
		7   => std_logic_vector(to_unsigned(0, 8)),
		8   => std_logic_vector(to_unsigned(0, 8)),
		9   => std_logic_vector(to_unsigned(0, 8)),
		10  => std_logic_vector(to_unsigned(0, 8)),
		11  => std_logic_vector(to_unsigned(0, 8)),
		12  => std_logic_vector(to_unsigned(0, 8)),
		13  => std_logic_vector(to_unsigned(0, 8)),
		14  => std_logic_vector(to_unsigned(0, 8)),
		15  => std_logic_vector(to_unsigned(0, 8)),
		16  => std_logic_vector(to_unsigned(0, 8)),
		17  => std_logic_vector(to_unsigned(0, 8)),
		18  => std_logic_vector(to_unsigned(0, 8)),
		19  => std_logic_vector(to_unsigned(0, 8)),
		20  => std_logic_vector(to_unsigned(0, 8)),
		21  => std_logic_vector(to_unsigned(0, 8)),
		22  => std_logic_vector(to_unsigned(1, 8)),
		23  => std_logic_vector(to_unsigned(1, 8)),
		24  => std_logic_vector(to_unsigned(1, 8)),
		25  => std_logic_vector(to_unsigned(1, 8)),
		26  => std_logic_vector(to_unsigned(1, 8)),
		27  => std_logic_vector(to_unsigned(1, 8)),
		28  => std_logic_vector(to_unsigned(1, 8)),
		29  => std_logic_vector(to_unsigned(2, 8)),
		30  => std_logic_vector(to_unsigned(2, 8)),
		31  => std_logic_vector(to_unsigned(2, 8)),
		32  => std_logic_vector(to_unsigned(2, 8)),
		33  => std_logic_vector(to_unsigned(2, 8)),
		34  => std_logic_vector(to_unsigned(2, 8)),
		35  => std_logic_vector(to_unsigned(3, 8)),
		36  => std_logic_vector(to_unsigned(3, 8)),
		37  => std_logic_vector(to_unsigned(3, 8)),
		38  => std_logic_vector(to_unsigned(3, 8)),
		39  => std_logic_vector(to_unsigned(3, 8)),
		40  => std_logic_vector(to_unsigned(4, 8)),
		41  => std_logic_vector(to_unsigned(4, 8)),
		42  => std_logic_vector(to_unsigned(4, 8)),
		43  => std_logic_vector(to_unsigned(4, 8)),
		44  => std_logic_vector(to_unsigned(5, 8)),
		45  => std_logic_vector(to_unsigned(5, 8)),
		46  => std_logic_vector(to_unsigned(5, 8)),
		47  => std_logic_vector(to_unsigned(5, 8)),
		48  => std_logic_vector(to_unsigned(6, 8)),
		49  => std_logic_vector(to_unsigned(6, 8)),
		50  => std_logic_vector(to_unsigned(6, 8)),
		51  => std_logic_vector(to_unsigned(7, 8)),
		52  => std_logic_vector(to_unsigned(7, 8)),
		53  => std_logic_vector(to_unsigned(7, 8)),
		54  => std_logic_vector(to_unsigned(8, 8)),
		55  => std_logic_vector(to_unsigned(8, 8)),
		56  => std_logic_vector(to_unsigned(8, 8)),
		57  => std_logic_vector(to_unsigned(9, 8)),
		58  => std_logic_vector(to_unsigned(9, 8)),
		59  => std_logic_vector(to_unsigned(9, 8)),
		60  => std_logic_vector(to_unsigned(10, 8)),
		61  => std_logic_vector(to_unsigned(10, 8)),
		62  => std_logic_vector(to_unsigned(11, 8)),
		63  => std_logic_vector(to_unsigned(11, 8)),
		64  => std_logic_vector(to_unsigned(11, 8)),
		65  => std_logic_vector(to_unsigned(12, 8)),
		66  => std_logic_vector(to_unsigned(12, 8)),
		67  => std_logic_vector(to_unsigned(13, 8)),
		68  => std_logic_vector(to_unsigned(13, 8)),
		69  => std_logic_vector(to_unsigned(13, 8)),
		70  => std_logic_vector(to_unsigned(14, 8)),
		71  => std_logic_vector(to_unsigned(14, 8)),
		72  => std_logic_vector(to_unsigned(15, 8)),
		73  => std_logic_vector(to_unsigned(15, 8)),
		74  => std_logic_vector(to_unsigned(16, 8)),
		75  => std_logic_vector(to_unsigned(16, 8)),
		76  => std_logic_vector(to_unsigned(17, 8)),
		77  => std_logic_vector(to_unsigned(17, 8)),
		78  => std_logic_vector(to_unsigned(18, 8)),
		79  => std_logic_vector(to_unsigned(18, 8)),
		80  => std_logic_vector(to_unsigned(19, 8)),
		81  => std_logic_vector(to_unsigned(19, 8)),
		82  => std_logic_vector(to_unsigned(20, 8)),
		83  => std_logic_vector(to_unsigned(21, 8)),
		84  => std_logic_vector(to_unsigned(21, 8)),
		85  => std_logic_vector(to_unsigned(22, 8)),
		86  => std_logic_vector(to_unsigned(22, 8)),
		87  => std_logic_vector(to_unsigned(23, 8)),
		88  => std_logic_vector(to_unsigned(23, 8)),
		89  => std_logic_vector(to_unsigned(24, 8)),
		90  => std_logic_vector(to_unsigned(25, 8)),
		91  => std_logic_vector(to_unsigned(25, 8)),
		92  => std_logic_vector(to_unsigned(26, 8)),
		93  => std_logic_vector(to_unsigned(27, 8)),
		94  => std_logic_vector(to_unsigned(27, 8)),
		95  => std_logic_vector(to_unsigned(28, 8)),
		96  => std_logic_vector(to_unsigned(29, 8)),
		97  => std_logic_vector(to_unsigned(29, 8)),
		98  => std_logic_vector(to_unsigned(30, 8)),
		99  => std_logic_vector(to_unsigned(31, 8)),
		100 => std_logic_vector(to_unsigned(31, 8)),
		101 => std_logic_vector(to_unsigned(32, 8)),
		102 => std_logic_vector(to_unsigned(33, 8)),
		103 => std_logic_vector(to_unsigned(34, 8)),
		104 => std_logic_vector(to_unsigned(34, 8)),
		105 => std_logic_vector(to_unsigned(35, 8)),
		106 => std_logic_vector(to_unsigned(36, 8)),
		107 => std_logic_vector(to_unsigned(37, 8)),
		108 => std_logic_vector(to_unsigned(37, 8)),
		109 => std_logic_vector(to_unsigned(38, 8)),
		110 => std_logic_vector(to_unsigned(39, 8)),
		111 => std_logic_vector(to_unsigned(40, 8)),
		112 => std_logic_vector(to_unsigned(40, 8)),
		113 => std_logic_vector(to_unsigned(41, 8)),
		114 => std_logic_vector(to_unsigned(42, 8)),
		115 => std_logic_vector(to_unsigned(43, 8)),
		116 => std_logic_vector(to_unsigned(44, 8)),
		117 => std_logic_vector(to_unsigned(45, 8)),
		118 => std_logic_vector(to_unsigned(46, 8)),
		119 => std_logic_vector(to_unsigned(46, 8)),
		120 => std_logic_vector(to_unsigned(47, 8)),
		121 => std_logic_vector(to_unsigned(48, 8)),
		122 => std_logic_vector(to_unsigned(49, 8)),
		123 => std_logic_vector(to_unsigned(50, 8)),
		124 => std_logic_vector(to_unsigned(51, 8)),
		125 => std_logic_vector(to_unsigned(52, 8)),
		126 => std_logic_vector(to_unsigned(53, 8)),
		127 => std_logic_vector(to_unsigned(54, 8)),
		128 => std_logic_vector(to_unsigned(55, 8)),
		129 => std_logic_vector(to_unsigned(56, 8)),
		130 => std_logic_vector(to_unsigned(57, 8)),
		131 => std_logic_vector(to_unsigned(58, 8)),
		132 => std_logic_vector(to_unsigned(59, 8)),
		133 => std_logic_vector(to_unsigned(60, 8)),
		134 => std_logic_vector(to_unsigned(61, 8)),
		135 => std_logic_vector(to_unsigned(62, 8)),
		136 => std_logic_vector(to_unsigned(63, 8)),
		137 => std_logic_vector(to_unsigned(64, 8)),
		138 => std_logic_vector(to_unsigned(65, 8)),
		139 => std_logic_vector(to_unsigned(66, 8)),
		140 => std_logic_vector(to_unsigned(67, 8)),
		141 => std_logic_vector(to_unsigned(68, 8)),
		142 => std_logic_vector(to_unsigned(69, 8)),
		143 => std_logic_vector(to_unsigned(70, 8)),
		144 => std_logic_vector(to_unsigned(71, 8)),
		145 => std_logic_vector(to_unsigned(72, 8)),
		146 => std_logic_vector(to_unsigned(73, 8)),
		147 => std_logic_vector(to_unsigned(74, 8)),
		148 => std_logic_vector(to_unsigned(76, 8)),
		149 => std_logic_vector(to_unsigned(77, 8)),
		150 => std_logic_vector(to_unsigned(78, 8)),
		151 => std_logic_vector(to_unsigned(79, 8)),
		152 => std_logic_vector(to_unsigned(80, 8)),
		153 => std_logic_vector(to_unsigned(81, 8)),
		154 => std_logic_vector(to_unsigned(83, 8)),
		155 => std_logic_vector(to_unsigned(84, 8)),
		156 => std_logic_vector(to_unsigned(85, 8)),
		157 => std_logic_vector(to_unsigned(86, 8)),
		158 => std_logic_vector(to_unsigned(88, 8)),
		159 => std_logic_vector(to_unsigned(89, 8)),
		160 => std_logic_vector(to_unsigned(90, 8)),
		161 => std_logic_vector(to_unsigned(91, 8)),
		162 => std_logic_vector(to_unsigned(93, 8)),
		163 => std_logic_vector(to_unsigned(94, 8)),
		164 => std_logic_vector(to_unsigned(95, 8)),
		165 => std_logic_vector(to_unsigned(96, 8)),
		166 => std_logic_vector(to_unsigned(98, 8)),
		167 => std_logic_vector(to_unsigned(99, 8)),
		168 => std_logic_vector(to_unsigned(100, 8)),
		169 => std_logic_vector(to_unsigned(102, 8)),
		170 => std_logic_vector(to_unsigned(103, 8)),
		171 => std_logic_vector(to_unsigned(104, 8)),
		172 => std_logic_vector(to_unsigned(106, 8)),
		173 => std_logic_vector(to_unsigned(107, 8)),
		174 => std_logic_vector(to_unsigned(109, 8)),
		175 => std_logic_vector(to_unsigned(110, 8)),
		176 => std_logic_vector(to_unsigned(111, 8)),
		177 => std_logic_vector(to_unsigned(113, 8)),
		178 => std_logic_vector(to_unsigned(114, 8)),
		179 => std_logic_vector(to_unsigned(116, 8)),
		180 => std_logic_vector(to_unsigned(117, 8)),
		181 => std_logic_vector(to_unsigned(119, 8)),
		182 => std_logic_vector(to_unsigned(120, 8)),
		183 => std_logic_vector(to_unsigned(121, 8)),
		184 => std_logic_vector(to_unsigned(123, 8)),
		185 => std_logic_vector(to_unsigned(124, 8)),
		186 => std_logic_vector(to_unsigned(126, 8)),
		187 => std_logic_vector(to_unsigned(128, 8)),
		188 => std_logic_vector(to_unsigned(129, 8)),
		189 => std_logic_vector(to_unsigned(131, 8)),
		190 => std_logic_vector(to_unsigned(132, 8)),
		191 => std_logic_vector(to_unsigned(134, 8)),
		192 => std_logic_vector(to_unsigned(135, 8)),
		193 => std_logic_vector(to_unsigned(137, 8)),
		194 => std_logic_vector(to_unsigned(138, 8)),
		195 => std_logic_vector(to_unsigned(140, 8)),
		196 => std_logic_vector(to_unsigned(142, 8)),
		197 => std_logic_vector(to_unsigned(143, 8)),
		198 => std_logic_vector(to_unsigned(145, 8)),
		199 => std_logic_vector(to_unsigned(146, 8)),
		200 => std_logic_vector(to_unsigned(148, 8)),
		201 => std_logic_vector(to_unsigned(150, 8)),
		202 => std_logic_vector(to_unsigned(151, 8)),
		203 => std_logic_vector(to_unsigned(153, 8)),
		204 => std_logic_vector(to_unsigned(155, 8)),
		205 => std_logic_vector(to_unsigned(157, 8)),
		206 => std_logic_vector(to_unsigned(158, 8)),
		207 => std_logic_vector(to_unsigned(160, 8)),
		208 => std_logic_vector(to_unsigned(162, 8)),
		209 => std_logic_vector(to_unsigned(163, 8)),
		210 => std_logic_vector(to_unsigned(165, 8)),
		211 => std_logic_vector(to_unsigned(167, 8)),
		212 => std_logic_vector(to_unsigned(169, 8)),
		213 => std_logic_vector(to_unsigned(170, 8)),
		214 => std_logic_vector(to_unsigned(172, 8)),
		215 => std_logic_vector(to_unsigned(174, 8)),
		216 => std_logic_vector(to_unsigned(176, 8)),
		217 => std_logic_vector(to_unsigned(178, 8)),
		218 => std_logic_vector(to_unsigned(179, 8)),
		219 => std_logic_vector(to_unsigned(181, 8)),
		220 => std_logic_vector(to_unsigned(183, 8)),
		221 => std_logic_vector(to_unsigned(185, 8)),
		222 => std_logic_vector(to_unsigned(187, 8)),
		223 => std_logic_vector(to_unsigned(189, 8)),
		224 => std_logic_vector(to_unsigned(191, 8)),
		225 => std_logic_vector(to_unsigned(193, 8)),
		226 => std_logic_vector(to_unsigned(194, 8)),
		227 => std_logic_vector(to_unsigned(196, 8)),
		228 => std_logic_vector(to_unsigned(198, 8)),
		229 => std_logic_vector(to_unsigned(200, 8)),
		230 => std_logic_vector(to_unsigned(202, 8)),
		231 => std_logic_vector(to_unsigned(204, 8)),
		232 => std_logic_vector(to_unsigned(206, 8)),
		233 => std_logic_vector(to_unsigned(208, 8)),
		234 => std_logic_vector(to_unsigned(210, 8)),
		235 => std_logic_vector(to_unsigned(212, 8)),
		236 => std_logic_vector(to_unsigned(214, 8)),
		237 => std_logic_vector(to_unsigned(216, 8)),
		238 => std_logic_vector(to_unsigned(218, 8)),
		239 => std_logic_vector(to_unsigned(220, 8)),
		240 => std_logic_vector(to_unsigned(222, 8)),
		241 => std_logic_vector(to_unsigned(224, 8)),
		242 => std_logic_vector(to_unsigned(227, 8)),
		243 => std_logic_vector(to_unsigned(229, 8)),
		244 => std_logic_vector(to_unsigned(231, 8)),
		245 => std_logic_vector(to_unsigned(233, 8)),
		246 => std_logic_vector(to_unsigned(235, 8)),
		247 => std_logic_vector(to_unsigned(237, 8)),
		248 => std_logic_vector(to_unsigned(239, 8)),
		249 => std_logic_vector(to_unsigned(241, 8)),
		250 => std_logic_vector(to_unsigned(244, 8)),
		251 => std_logic_vector(to_unsigned(246, 8)),
		252 => std_logic_vector(to_unsigned(248, 8)),
		253 => std_logic_vector(to_unsigned(250, 8)),
		254 => std_logic_vector(to_unsigned(252, 8)),
		255 => std_logic_vector(to_unsigned(255, 8))
	);
begin
	pixelData_out  <= gamma_table(to_integer(unsigned(pixelData_in)));
end architecture RTL;
